`include "svlib_private_base_pkg.sv"
`include "svlib_pkg_Str.sv"
`include "svlib_pkg_Regex.sv"
`include "svlib_pkg_Enum.sv"
`include "svlib_pkg_File.sv"
`include "svlib_pkg_Sys.sv"
`include "svlib_pkg_Cfg.sv"
