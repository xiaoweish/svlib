`ifndef SVLIB_MACROS__DEFINED
`define SVLIB_MACROS__DEFINED

`define forenum(E,e,i=foreach_enum_position_iterator) \
  for (E e = e.first, int i=0; i<e.num; e=e.next, i++)
  
`define SVLIB_CLASS(T, B)                         \
  class T extends B;                              \
    protected static function T randstable_new(); \
      `ifdef SVLIB_NO_RANDSTABLE_NEW              \
      T result = new();                           \
      `else                                       \
      std::process p = std::process::self();      \
      string randstate = p.get_randstate();       \
      T result = new();                           \
      p.set_randstate(randstate);                 \
      `endif                                      \
      return result;                              \
    endfunction                                   \

`endif
