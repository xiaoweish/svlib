`ifndef SVLIB_STR_PKG__DEFINED
`define SVLIB_STR_PKG__DEFINED

`define SVLIB_NO_RANDSTABLE_NEW

`include "svlib_macros.sv"

package svlib_Str_pkg;

  import "DPI-C" function int SvLib_regexRun(
                           input  string re,
                           input  string str,
                           input  int    cflags,
                           input  int    startPos,
                           output int    matchCount,
                           output int    matchList[]);
  import "DPI-C" function string SvLib_regexErrorString(input int err);

  typedef string qs[$];
  
  function automatic bit isspace(byte unsigned ch);
    return (ch inside {"\t", "\n", "\r", " ", 160});  // nbsp
  endfunction
  
  virtual class svlib_base;// #(parameter type T = int);
    /*protected T*/ svlib_base obstack_link;
    /*
    protected static function T randstable_new();
      `ifdef SVLIB_NO_RANDSTABLE_NEW
      T result = new();
      `else
      std::process p = std::process::self();
      string randstate = p.get_randstate();
      T result = new();
      p.set_randstate(randstate);
      `endif
      return result;
    endfunction
    */
  endclass
  
  virtual class Obstack #(parameter type T=int);
    local static svlib_base head;//T   head;
    local static int constructed_ = 0;
    local static int get_calls_ = 0;
    local static int put_calls_ = 0;
    
    static function T get();
      T result;
      if (head == null) begin
        result = T::create();
        constructed_++;
      end
      else begin
        $cast(result, head);//result = head;
        head = head.obstack_link;
      end
      get_calls_++;
      return result;
    endfunction
    static function void put(T t);
      put_calls_++;
      if (t == null) return;
      t.obstack_link = head;
      head = t;
    endfunction
    // debug/test only - DO NOT USE normally
    static function void stats(
        output int depth,
        output int constructed,
        output int get_calls,
        output int put_calls
      );
      /*T*/svlib_base p = head;
      depth = 0;
      while (p != null) begin
        depth++;
        p = p.obstack_link;
      end
      constructed = constructed_;
      get_calls = get_calls_;
      put_calls = put_calls_;
    endfunction
  endclass
  
  // Str: various string manipulations.
  // Most functions come in two flavors:
  // - a package version named str_XXX that takes a string value,
  //   does some work on it and returns a result; and
  // - an object version named .XXX that operates on a stored
  //   Str object, possibly returning a result and possibly
  //   modifying the stored object.
  //
  typedef class Str;
  class Str extends svlib_base;//#(Str);
  
    typedef enum {NONE, LEFT, RIGHT, BOTH} side_e;
    typedef enum {START, END} origin_e;
  
    // Save a string as an object so that further manipulations can
    // be performed on it.  Get and set the object's string value.
    extern static  function Str    create(string s = "");
    extern virtual function string get();
    extern virtual function Str    copy();
    extern virtual function int    len();
    
    extern virtual function void   set(string s);
    
    extern virtual function void   append(string s);

    // Find the first occurrence of substr in s, starting from the "start"
    // position. If a match is found, return the index of the first character
    // of the match.  If no match is found, return -1.
    extern virtual function int    first(string substr, int ignore=0);
    extern virtual function int    last (string substr, int ignore=0);
    
    // Split a string on every occurrence of a given character
    extern virtual function qs     split(string splitset="", bit keepSplitters=0);
    
    // Get a range (substring). The starting position 'p' is an anchor point,
    // like an I-beam cursor, just to the left of the specified character.
    // If 'origin' is START, count 'p' from the left end of the string, 
    // with its value increasing towards the right. If 'origin' is END, 
    // count 'p' from the right end of the string, with its value increasing
    // towards the left.
    // The range size 'n' specifies a count of characters to the right of 'p',
    // or to the left of 'p' if 'n' is negative; n==0 specifies an empty string.
    // If p<0, treat it as the corresponding number of character positions
    // beyond the end (or start) of the string.
    // Clip result to smaller than n if necessary so that the result remains
    // entirely within the bounds of the original string.
    extern virtual function string range(int p, int n, origin_e origin=START);
    
    // Replace the range p/n with some other string, not necessarily same length.
    // If n==0 this is an insert operation.
    extern virtual function void   replace(string rs, int p, int n, origin_e origin=START);
    
    // Tokenize a string on whitespace boundaries
    extern virtual function qs     tokens();
    
    // Trim a string (remove leading and/or trailing whitespace)
    extern virtual function void   trim(side_e side=BOTH);
    
    // Justify a string (pad to width with spaces on left/right/both)
    extern virtual function void   just(int width, side_e side=BOTH);
    
    protected string value;
    
    extern protected function void get_range_positions(
      int p, int n, origin_e origin=START,
      output int L, output int R
    );
    extern protected function void clip_to_bounds(inout int n);
    
  endclass
  
  typedef class Regex;
  class Regex extends svlib_base;//#(Regex);
  
    extern static  function Regex  create(string s = "", bit nocase=0, bit noline=0);
    extern virtual function void   setRE(string s);
    extern virtual function void   setOpts(bit nocase, bit noline);
//    extern virtual function void   setMaxMatches(int maxMatches);
    
    extern virtual function string getRE();
    extern virtual function void   getOpts(output bit nocase, output bit noline);
//    extern virtual function int    getMaxMatches();
    extern virtual function Regex  copy();
    
    extern virtual function void   purge();
    
    extern virtual function int    run(Str s, output int nMatches, input int startPos=0);
    extern virtual function int    getMatchPosition(int match, output int L, output int R);
    extern virtual function int    getMatchString(int match, output string s);
    extern virtual function string getErrorString();
    
    protected int lastMatchCount;
    protected int lastError;
    protected int matchList[20];
    protected Str runStr;
    
    protected int     compiledRegexKey;    // for lookup on C side
    protected chandle compiledRegexHandle; // check on C-side pointer
    
    protected bit    nocase;
    protected bit    noline;
    protected string text;
  
  endclass

  
  function void Str::get_range_positions(
    int p, int n, origin_e origin=START,
    output int L, output int R
  );
    int len = value.len;
    // establish start position "just to the left of"
    if (origin==END) begin
      L = len - p;
    end
    else begin
      L = p;
    end
    // establish L/R boundaries
    R = L;
    if (n<0) begin
      // 'p' is right end, push L leftwards appropriately
      L += n;
    end
    else begin
      // 'p' is left end, push R rightwards appropriately
      R += n;
    end
  endfunction

  function void Str::clip_to_bounds(inout int n);
    if (n<0) n=0; else if (n>value.len) n=value.len;
  endfunction

  // Save a string as an object so that further manipulations can
  // be performed on it.
  function Str Str::create(string s = "");
    Str result = new;//randstable_new();
    result.set(s);
    return result;
  endfunction

  // Get the object's string value.
  function string Str::get();
    return value;
  endfunction

  // Get the string's length.
  function int Str::len();
    return value.len;
  endfunction
  
  function Str Str::copy(); 
    return create(value);
  endfunction

  function void Str::set(string s);
    value = s;
  endfunction

  function void Str::append(string s);
    replace(s, 0, 0, END);
  endfunction


  // Find the first occurrence of substr in s, starting from the "start"
  // position. If a match is found, return the index of the first character
  // of the match.  If no match is found, return -1.
  function int Str::first(string substr, int ignore=0);
    for (int i=ignore; i<=(value.len-substr.len); i++) begin
      if (substr == value.substr(i, i+substr.len-1)) return i;
    end
    return -1;
  endfunction

  function int Str::last(string substr, int ignore=0);
    for (int i=(value.len-substr.len)-ignore; i>=0; i--) begin
      if (substr == value.substr(i, i+substr.len-1)) return i;
    end
    return -1;
  endfunction

  // Replace the range p/n with some other string, not necessarily same length
  function void Str::replace(string rs, int p, int n, origin_e origin=START);
    int len = value.len;
    int L, R;
    get_range_positions(p, n, origin, L, R);
    clip_to_bounds(L);
    clip_to_bounds(R);
    value = {value.substr(0, L-1), rs, value.substr(R, len-1)};
  endfunction
  //
  function automatic string str_replace(
      string orig, string rs, int p, int n=0, Str::origin_e origin=Str::START
    );
    Str obj = Obstack#(Str)::get();
    obj.set(orig);
    obj.replace(rs, p, n, origin);
    str_replace = obj.get();
    Obstack#(Str)::put(obj);
  endfunction

  function string Str::range(int p, int n, origin_e origin=START);
    int L, R;
    get_range_positions(p, n, origin, L, R);
    clip_to_bounds(L);
    clip_to_bounds(R);
    // adjust for substr conventions
    R--;
    return value.substr(L, R);
  endfunction

  // Trim a string (remove leading and/or trailing whitespace)
  function void Str::trim(side_e side=BOTH);
    int first;
    int last;
    if (side == NONE) return;
    first = 0;
    last  = value.len-1;
    if (side inside {LEFT, BOTH}) begin
      while ((first <= last) && isspace(value[first])) first++;
    end
    if (side inside {RIGHT, BOTH}) begin
      while ((first <= last) && isspace(value[last])) last--;
    end
    value = value.substr(first, last);
  endfunction

  // Justify a string (pad to width with spaces on left/right/both)
  function void Str::just(int width, side_e side=BOTH);
    int n, n2;
    if (side == NONE) return;
    n = width - signed'(value.len);
    if (n <= 0) return;
    case (side)
      RIGHT:
        value = { {n{" "}}, value };
      LEFT:
        value = { value, {n{" "}} };
      BOTH:
        begin
          n2 = n/2;
          value = { {n2{" "}}, value, {n-n/2{" "}} };
        end
    endcase
  endfunction
    
  // Split a string on every occurrence of a given character
  function qs Str::split(string splitset="", bit keepSplitters=0);
    split = {};
    if (splitset == "") begin
      for (int i=0; i<value.len(); i++) begin
        split.push_back(value.substr(i,i));
      end
    end
    else begin
      byte unsigned splitchars[$];
      int anchor = 0;
      foreach (splitset[i]) begin
        splitchars.push_back(splitset[i]);
      end
      foreach (value[i]) begin
        if (value[i] inside {splitchars}) begin
          split.push_back(value.substr(anchor, i-1));
          if (keepSplitters) begin
            split.push_back(value.substr(i,i));
          end
          anchor = i+1;
        end
      end
      split.push_back(value.substr(anchor, value.len()-1));
    end
  endfunction


  function Regex  Regex::create(string s = "", bit nocase=0, bit noline=0);
    Regex r = new(); //randstable_new();
    r.setRE(s);
    r.setOpts(nocase, noline);
//    r.setMaxMatches(10);  // sensible default
    return r;
  endfunction
  
  function void   Regex::setRE(string s);
    if (s!=text) begin
      // RE text has changed, so we must reset the object
      this.text = s;
      purge();
    end
  endfunction
  
  function void   Regex::setOpts(bit nocase, bit noline);
    if (nocase!=nocase || noline!=noline) begin
      // Something has changed, so we must reset the object
      this.nocase = nocase;
      this.noline = noline;
      purge();
    end
  endfunction
  
//   function void   Regex::setMaxMatches(int maxMatches);
//     if (maxMatches*2 != matchList.size()) begin
//       matchList = new[maxMatches*2];
//     end
//   endfunction
  
  function void   Regex::purge();
    compiledRegexHandle = null;
    lastMatchCount = -1; // Not matched at all
    lastError = -1;  // No match attempt
  endfunction
  
  function string Regex::getRE();
    return text;
  endfunction
  
  function void   Regex::getOpts(output bit nocase, output bit noline);
    nocase = this.nocase;
    noline = this.noline;
  endfunction
  
//   function int    Regex::getMaxMatches();
//     return matchList.size()/2;
//   endfunction
  
  function Regex  Regex::copy();
    Regex it = create(text, nocase, noline);
//    it.setMaxMatches(getMaxMatches());
  endfunction
  
  // REVISIT Incomplete implementations:
  
  // Tokenize a string on whitespace boundaries. Commas and
  // string quotes are respected, CSV-fashion.
  function qs Str::tokens();
    return {};
  endfunction
  
  function int    Regex::run(Str s, output int nMatches, input int startPos=0);
    int result;
    runStr = s;
    nMatches = 0;
    lastMatchCount = -1;  // pessimistic
    
    lastError = SvLib_regexRun(
      .re(text), .str(s.get()), .cflags(0), .startPos(startPos), 
      .matchCount(nMatches), .matchList(matchList));
    for (int i=2*nMatches; i<$size(matchList,1); i++) matchList[i] = -1;
    
    $display("result from Regex::run = %0d, nMatches=%0d", lastError, nMatches);
    if (lastError) return lastError;
    
    for (int i=0; i<$size(matchList,1); i+=2) begin
      $display("match %0d - %0d:%0d", i/2, matchList[i], matchList[i+1]);
    end
    lastMatchCount = nMatches;
    return 0;
  endfunction
  
  function int    Regex::getMatchPosition(int match, output int L, output int R);
    if (match>lastMatchCount || match<0) begin
      L = -1;
      R = -1;
      return 1;
    end
    else begin
      L = matchList[match*2];
      R = matchList[match*2+1] - 1;
      return 0;
    end
  endfunction
  
  function int    Regex::getMatchString(int match, output string s);
    int L, R, result;
    s = "";
    result = getMatchPosition(match, L, R);
    if (result) return result;
    if (runStr == null) return 1;
    s = runStr.range(L, R+1-L);
    return 0;
  endfunction
  
  function string Regex::getErrorString();
    case (lastError)
      0  : return "";
      -1 : return "SvLib_regex not yet run";
      default :
        return SvLib_regexErrorString(lastError);
    endcase
  endfunction
    
endpackage

`endif
